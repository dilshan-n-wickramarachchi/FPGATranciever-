module receiver#(
			//Local Parameters 
			parameter RX_STATE_START	= 2'b00,
			parameter RX_STATE_DATA		= 2'b01,
			parameter RX_STATE_STOP		= 2'b10
		)(
		//Input Wires 
		input wire rx,
		input wire rdy_clr,
		input wire clk_50m,
		input wire clken,
		//Ouput registers 
		output reg rdy,
		output reg [7:0] data);

initial begin
	rdy = 0;
	data = 8'b0;
end



reg [1:0] state = RX_STATE_START;
reg [3:0] sample = 0;
reg [3:0] bitpos = 0;
reg [7:0] scratch = 8'b0;

always @(posedge clk_50m) begin
	if(rdy_clr)begin
		rdy<=0;
		if (clken) begin
			case (state)
			RX_STATE_START: begin
				/*
				* Start counting from the first low sample, once we've
				* sampled a full bit, start collecting data bits.
				*/
				if (!rx || sample != 0)
					sample <= sample + 4'b1;

				if (sample == 15) begin
					state <= RX_STATE_DATA;
					bitpos <= 0;
					sample <= 0;
					scratch <= 0;
				end
			end
			RX_STATE_DATA: begin
				sample <= sample + 4'b1;
				if (sample == 4'h8) begin
					scratch[bitpos[2:0]] <= rx;
					bitpos <= bitpos + 4'b1;
				end
				if (bitpos == 8 && sample == 15)
					state <= RX_STATE_STOP;
			end
			RX_STATE_STOP: begin
				/*
				 * Our baud clock may not be running at exactly the
				 * same rate as the transmitter.  If we thing that
				 * we're at least half way into the stop bit, allow
				 * transition into handling the next start bit.
				 */
				if (sample == 15 || (sample >= 8 && !rx)) begin
					state <= RX_STATE_START;
					data <= scratch; 
					sample <= 0;
				end else begin
					sample <= sample + 4'b1;
				end
			end
			default: begin
				state <= RX_STATE_START;
			end
			endcase
		end 
		
	end else begin
		rdy<=1;
		data = 8'b0;
	end
end
endmodule

